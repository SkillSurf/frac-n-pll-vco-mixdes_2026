** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/top-pll/LCVCO_DSM_tb.sch
**.subckt LCVCO_DSM_tb OUTn VDD VCTRL GND Ibias
*.opin OUTn
*.iopin VDD
*.iopin VCTRL
*.iopin GND
*.iopin Ibias
V1 VDD GND 1.2
V2 VCTRL GND pulse(0.3 1.0 50n 100n 100n 200n)
I0 VDD Ibias 50u
x5 OUTp net7 VDD GND sg13g2_inv_2
x1 VDD net7 OUTn Ibias VCTRL GND LC_VCO
adut [ net1 net2 net3 net4 net5 ] [ net6 ] null dut
.model dut d_cosim simulation=./../dsm_and_freq_divider.so
A1 [ OUTp ] [ net1 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=0.6
A2 [ rst ] [ net2 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=0.6
A3 [ sclk ] [ net3 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=0.6
A4 [ sdata ] [ net4 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=0.6
A5 [ en ] [ net5 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=0.6
A6 [ net6 ] [ outd ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
* noconn rst
* noconn sclk
* noconn sdata
* noconn en
**** begin user architecture code



.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ_stat
.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice
.global VDD GND






.include ./IHP_4nH_Inductor.spice
.param temp=27
.save v(OUTp) v(Vctrl)
.save v(dout) v(sdata) v(sclk) v(en) v(rst)
.save v(dsm_clk) v(outd)
.control
.options maxstep=50p reltol=1e-3 abstol=1e-6

*.ic v(OUTp)=0.6
tran 0.5n 1m
remzerovec
linearize v(OUTp) v(Vctrl) v(outd)

    let n_pts = length(time)
    let freq_vector = unitvec(n_pts) * 0

    * Advanced script to calculate instantaneous frequency
    let i = 1
    let last_cross = 0
    while i < length(time)
        if (v(OUTp)[i] >= 0.6) & (v(OUTp)[i-1] < 0.6)
            let current_cross = time[i]
            let period = current_cross - last_cross
            let inst_freq = 1 / period
            let freq_vector[i] = inst_freq
            let last_cross = current_cross
        else
            let freq_vector[i] = freq_vector[i-1]
        end
        let i = i + 1
    end

* Save transient waveform to raw file
write LCVCO_DSM.raw

*quit 0
.endc


* to generate following file copy stimuli.test
* to the simulation directory and run simulation -> Utile Stimuli Editor (GUI),
* and press 'Translate'
.include stimuli_test.cir


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/lc-vco/LC_VCO.sym # of pins=6
** sym_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/lc-vco/LC_VCO.sym
** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/lc-vco/LC_VCO.sch
.subckt LC_VCO VDD OUTp OUTn Ibias VCTRL GND
*.iopin VDD
*.opin OUTp
*.opin OUTn
*.iopin GND
*.iopin VCTRL
*.iopin Ibias
XM6 net1 Ibias GND GND sg13_lv_nmos w=1u l=0.15u ng=1 m=60
XM5 Ibias Ibias GND GND sg13_lv_nmos w=1u l=0.15u ng=1 m=1
XM4 OUTp OUTn VDD VDD sg13_lv_pmos w=8.5u l=0.5u ng=1 m=13
X5M3 OUTn OUTp VDD VDD sg13_lv_pmos w=8.5u l=0.5u ng=1 m=13
XM2 OUTp OUTn net1 GND sg13_lv_nmos w=2u l=0.5u ng=1 m=12
XM1 OUTn OUTp net1 GND sg13_lv_nmos w=2u l=0.5u ng=1 m=12
XC3 OUTp OUTn cap_cmim w=4.0e-6 l=4.0e-6 m=13.6
XMv2 OUTp VCTRL OUTp VDD sg13_lv_pmos w=4u l=4u ng=1 m=22
XMv1 OUTn VCTRL OUTn VDD sg13_lv_pmos w=4u l=4u ng=1 m=22
*  x1 -  ihp_4nh_inductor  IS MISSING !!!!
XR1 OUTn OUTp sub! rhigh w=1e-6 l=1e-6 m=1.23 b=0
.ends

.GLOBAL GND
.GLOBAL VDD
.GLOBAL VCTRL
.GLOBAL Ibias
.end
