** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/lc-vco/LC_VCO_tb.sch
**.subckt LC_VCO_tb OUTp OUTn VDD VCTRL GND Ibias
*.opin OUTp
*.opin OUTn
*.iopin VDD
*.iopin VCTRL
*.iopin GND
*.iopin Ibias
V1 VDD GND 1.2
V2 VCTRL GND 0.6
x1 VDD OUTp OUTn Ibias VCTRL GND LC_VCO
I0 VDD Ibias 50u
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt
.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ_stat



.include ./IHP_4nH_Inductor.spice
.param temp=27
.control
save all
.ic v(OUTp)=0.6

.options maxstep=10n reltol=1e-3 abstol=1e-6
save v(vout)
tran 0.01n 0.5u UIC

* Save transient waveform to raw file
write LC_VCO_tb.raw

* Plot time-domain waveform
plot v(OUTp) xlimit 5n 60n

* Perform FFT on output
fft v(OUTp)

* Convert FFT magnitude to dB
let vmag = db(mag(v(OUTp)))

* Plot FFT result
plot vmag xlabel 'Frequency (Hz)' xlimit 0 5G

* Save FFT data to text file
wrdata fft_output(VCTRL=0.6).txt vmag

.endc


**** end user architecture code
**.ends

* expanding   symbol:  LC_VCO.sym # of pins=6
** sym_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/lc-vco/LC_VCO.sym
** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/lc-vco/LC_VCO.sch
.subckt LC_VCO VDD OUTp OUTn Ibias VCTRL GND
*.iopin VDD
*.opin OUTp
*.opin OUTn
*.iopin GND
*.iopin VCTRL
*.iopin Ibias
XM6 net1 Ibias GND GND sg13_lv_nmos w=1u l=0.15u ng=1 m=60
XM5 Ibias Ibias GND GND sg13_lv_nmos w=1u l=0.15u ng=1 m=1
XM4 OUTp OUTn VDD VDD sg13_lv_pmos w=8.5u l=0.5u ng=1 m=13
X5M3 OUTn OUTp VDD VDD sg13_lv_pmos w=8.5u l=0.5u ng=1 m=13
XM7 OUTp OUTn net1 GND sg13_lv_nmos w=2u l=0.5u ng=1 m=12
XM8 OUTn OUTp net1 GND sg13_lv_nmos w=2u l=0.5u ng=1 m=12
XC3 OUTp OUTn cap_cmim w=4.0e-6 l=4.0e-6 m=10
R6 OUTp OUTn 1.25k m=1
R1 OUTp net2 4 m=1
x1 OUTn net2 ihp_4nh_inductor
XMv2 OUTp VCTRL OUTp VDD sg13_lv_pmos w=8u l=8u ng=1 m=35
XMv1 OUTn VCTRL OUTn VDD sg13_lv_pmos w=8u l=8u ng=1 m=35
.ends

.GLOBAL GND
.GLOBAL VDD
.GLOBAL VCTRL
.GLOBAL Ibias
.end
