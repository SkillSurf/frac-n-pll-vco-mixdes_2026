** sch_path: /foss/designs/iic-osic-tools/Analog_designs/LC-VCO-3Ghz/Design/design_data/xschem/LC_VCO_tb.sch
**.subckt LC_VCO_tb OUTp OUTn VDD VCTRL GND Ibias
*.opin OUTp
*.opin OUTn
*.iopin VDD
*.iopin VCTRL
*.iopin GND
*.iopin Ibias
V1 VDD GND 1.8
V2 VCTRL GND 0.9
x1 VDD OUTp OUTn Ibias VCTRL GND LC_VCO
I0 VDD Ibias 50u
**** begin user architecture code


.param temp=27
.options maxstep=10n reltol=1e-3 abstol=1e-6

.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.tran 0.01n 0.3u

* Save differential and single-ended outputs
.save v(OUTp) v(OUTn)

.control
  run
  * Save transient waveform to raw file
  write LC_VCO_tb.raw

  * Plot time-domain waveform
  plot v(OUTp) xlimit 0.0n 60n

  * Perform FFT on output
  fft v(OUTp)

  * Convert FFT magnitude to dB
  let vmag = db(mag(v(OUTp)))

  * Plot FFT result
  plot vmag xlabel 'Frequency (Hz)' xlimit 0 5G

  * Save FFT data to text file
  wrdata fft_output(VCTRL=0.9).txt vmag
.endc




**** end user architecture code
**.ends

* expanding   symbol:  LC_VCO.sym # of pins=6
** sym_path: /foss/designs/iic-osic-tools/Analog_designs/LC-VCO-3Ghz/Design/design_data/xschem/LC_VCO.sym
** sch_path: /foss/designs/iic-osic-tools/Analog_designs/LC-VCO-3Ghz/Design/design_data/xschem/LC_VCO.sch
.subckt LC_VCO VDD OUTp OUTn Ibias VCTRL GND
*.iopin VDD
*.opin OUTp
*.opin OUTn
*.iopin GND
*.iopin VCTRL
*.iopin Ibias
XM2 OUTn OUTp net1 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=18 m=18
XM3 OUTp OUTn net1 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=18 m=18
XM6 Ibias Ibias GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 net1 Ibias GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=60 m=60
L3 net2 OUTn 2n m=1
R5 OUTp net2 0.28 m=1
R6 OUTp OUTn 0.65k m=1
XC2 OUTp OUTn sky130_fd_pr__cap_mim_m3_2 W=4.5 L=4.5 MF=25 m=25
XM4 OUTp OUTn VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.74 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=21 m=21
XM1 OUTn OUTp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.74 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=21 m=21
XM5 OUTn VCTRL OUTn VDD sky130_fd_pr__pfet_01v8_lvt L=3 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=42 m=42
XC6 OUTn GND sky130_fd_pr__cap_mim_m3_2 W=1 L=1 MF=170 m=170
XM7 OUTp VCTRL OUTp VDD sky130_fd_pr__pfet_01v8_lvt L=3 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=42 m=42
XC1 OUTp GND sky130_fd_pr__cap_mim_m3_2 W=1 L=1 MF=170 m=170
.ends

.GLOBAL GND
.GLOBAL VDD
.GLOBAL VCTRL
.GLOBAL Ibias
.end
