** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/top-pll/PFD_CP_LCVCO_tb.sch
**.subckt PFD_CP_LCVCO_tb OUTn VDD VCTRL GND Ibias
*.opin OUTn
*.iopin VDD
*.iopin VCTRL
*.iopin GND
*.iopin Ibias
V1 VDD GND 1.2
V2 VCTRL GND pulse(0.3 1.0 50n 100n 100n 200n)
I0 VDD Ibias 50u
x5 OUTp net1 VDD GND sg13g2_inv_2
x1 VDD net1 OUTn Ibias VCTRL GND LC_VCO
x2 OUTp OUTd Freq_Div_std
**** begin user architecture code



.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ_stat
.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice
.global VDD GND






.model freq_div freq_div
.include ./IHP_4nH_Inductor.spice
.param temp=27
.control
pre_osdi ./freq_div.osdi
save all
*.ic v(OUTp)=0.6

tran 1p 200n UIC

linearize v(OUTp) v(Vctrl) v(outd)

    let n_pts = length(time)
    let freq_vector = unitvec(n_pts) * 0

    * Advanced script to calculate instantaneous frequency
    let i = 1
    let last_cross = 0
    while i < length(time)
        if (v(OUTp)[i] >= 0.6) & (v(OUTp)[i-1] < 0.6)
            let current_cross = time[i]
            let period = current_cross - last_cross
            let inst_freq = 1 / period
            let freq_vector[i] = inst_freq
            let last_cross = current_cross
        else
            let freq_vector[i] = freq_vector[i-1]
        end
        let i = i + 1
    end

* Save transient waveform to raw file
write LCVCO_freqdiv.raw

*quit 0
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/lc-vco/LC_VCO.sym # of pins=6
** sym_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/lc-vco/LC_VCO.sym
** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/lc-vco/LC_VCO.sch
.subckt LC_VCO VDD OUTp OUTn Ibias VCTRL GND
*.iopin VDD
*.opin OUTp
*.opin OUTn
*.iopin GND
*.iopin VCTRL
*.iopin Ibias
XM6 net1 Ibias GND GND sg13_lv_nmos w=1u l=0.15u ng=1 m=60
XM5 Ibias Ibias GND GND sg13_lv_nmos w=1u l=0.15u ng=1 m=1
XM4 OUTp OUTn VDD VDD sg13_lv_pmos w=8.5u l=0.5u ng=1 m=13
X5M3 OUTn OUTp VDD VDD sg13_lv_pmos w=8.5u l=0.5u ng=1 m=13
XM2 OUTp OUTn net1 GND sg13_lv_nmos w=2u l=0.5u ng=1 m=12
XM1 OUTn OUTp net1 GND sg13_lv_nmos w=2u l=0.5u ng=1 m=12
XC3 OUTp OUTn cap_cmim w=4.0e-6 l=4.0e-6 m=13.6
XMv2 OUTp VCTRL OUTp VDD sg13_lv_pmos w=4u l=4u ng=1 m=22
XMv1 OUTn VCTRL OUTn VDD sg13_lv_pmos w=4u l=4u ng=1 m=22
*  x1 -  ihp_4nh_inductor  IS MISSING !!!!
XR1 OUTn OUTp sub! rhigh w=1e-6 l=1e-6 m=1.23 b=0
.ends


* expanding   symbol:  /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/top-pll/FD/Freq_Div_std.sym # of
*+ pins=2
** sym_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/top-pll/FD/Freq_Div_std.sym
** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/top-pll/FD/Freq_Div_std.sch
.subckt Freq_Div_std F_IN F_OUT
*.opin F_OUT
*.ipin F_IN
x6 net3 net1 F_IN net1 VDD VDD GND sg13g2_dfrbp_1
x5 net4 net2 net3 net2 VDD VDD GND sg13g2_dfrbp_2
x7 net6 net5 net4 net5 VDD VDD GND sg13g2_dfrbp_2
x8 F_OUT net7 net6 net7 VDD VDD GND sg13g2_dfrbp_2
.ends

.GLOBAL GND
.GLOBAL VDD
.GLOBAL VCTRL
.GLOBAL Ibias
.end
