** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/top-pll/pll_temp_fredivider.sch
**.subckt pll_temp_fredivider OUTn
*.opin OUTn
V1 VDD GND 1.2
I0 VDD IbiasVCO 50u
Vfref F_REF GND 0 pulse(0 1.2 0n 0.1n 0.1n 5n 10n)
I1 Ibias GND 10m
R1 F_VCO F_DIV 4 m=1
x5 OUTp net1 VDD GND sg13g2_inv_2
x1 VDD net1 OUTn IbiasVCO CTRL GND LC_VCO
x2 VDD UP CTRL DN GND Ibias CP
x3 VDD UP F_REF F_VCO DN GND PFD_std
x4 OUTp F_DIV Freq_Div_std
**** begin user architecture code



.lib cornerMOSlv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ_stat
.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice
.global VDD GND


.param CP_N_L = 0.5u
.param CP_N_W = 60u
.param CP_P_M = 1
.param CP_P_L = 0.5u
.param CP_P_W = 200u
.param CP_N_M = 1
.param C_CP = 700p





.model freq_div freq_div
.include ./IHP_4nH_Inductor.spice
.option temp = 27
.param VDD = 1.2
.ic v(OUTp)=0.6

.control
.options maxstep=100P reltol=1e-3 abstol=1e-6
pre_osdi ./freq_div.osdi
save v(CTRL) v(OUTp) v(F_REF) v(F_DIV) v(UP) v(DN) v(F_VCO)

tran 50p 500n uic
write tb_pll_freq_div.raw
*quit 0
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/lc-vco/LC_VCO.sym # of pins=6
** sym_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/lc-vco/LC_VCO.sym
** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/lc-vco/LC_VCO.sch
.subckt LC_VCO VDD OUTp OUTn Ibias VCTRL GND
*.iopin VDD
*.opin OUTp
*.opin OUTn
*.iopin GND
*.iopin VCTRL
*.iopin Ibias
XM6 net1 Ibias GND GND sg13_lv_nmos w=1u l=0.15u ng=1 m=60
XM5 Ibias Ibias GND GND sg13_lv_nmos w=1u l=0.15u ng=1 m=1
XM4 OUTp OUTn VDD VDD sg13_lv_pmos w=8.5u l=0.5u ng=1 m=13
X5M3 OUTn OUTp VDD VDD sg13_lv_pmos w=8.5u l=0.5u ng=1 m=13
XM2 OUTp OUTn net1 GND sg13_lv_nmos w=2u l=0.5u ng=1 m=12
XM1 OUTn OUTp net1 GND sg13_lv_nmos w=2u l=0.5u ng=1 m=12
XC3 OUTp OUTn cap_cmim w=4.0e-6 l=4.0e-6 m=13.6
XMv2 OUTp VCTRL OUTp VDD sg13_lv_pmos w=4u l=4u ng=1 m=22
XMv1 OUTn VCTRL OUTn VDD sg13_lv_pmos w=4u l=4u ng=1 m=22
*  x1 -  ihp_4nh_inductor  IS MISSING !!!!
XR1 OUTn OUTp sub! rhigh w=1e-6 l=1e-6 m=1.23 b=0
.ends


* expanding   symbol:  /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/charge-pump/CP.sym # of pins=6
** sym_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/charge-pump/CP.sym
** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/charge-pump/CP.sch
.subckt CP VDD UP CTRL DN GND Ibias
*.opin CTRL
*.ipin UP
*.ipin VDD
*.ipin Ibias
*.ipin DN
*.ipin GND
XM2 Vbn Vbn net2 GND sg13_lv_nmos w={CP_N_W} l={CP_N_L} ng=1 m={CP_N_M}
XM1 net2 VDD GND GND sg13_lv_nmos w={CP_N_W} l={CP_N_L} ng=1 m={CP_N_M}
XM3 Vbn Vbp net1 VDD sg13_lv_pmos w={CP_P_W} l={CP_P_L} ng=1 m={CP_P_M}
XM4 net1 GND VDD VDD sg13_lv_pmos w={CP_P_W} l={CP_P_L} ng=1 m={CP_P_M}
XM7 Vbp Vbp net7 VDD sg13_lv_pmos w={CP_P_W} l={CP_P_L} ng=1 m={CP_P_M}
XM8 net7 GND VDD VDD sg13_lv_pmos w={CP_P_W} l={CP_P_L} ng=1 m={CP_P_M}
XM5 net6 Vbn net3 GND sg13_lv_nmos w={CP_N_W} l={CP_N_L} ng=1 m={CP_N_M}
XM6 net3 DN GND GND sg13_lv_nmos w={CP_N_W} l={CP_N_L} ng=1 m={CP_N_M}
XM9 net6 Vbp net4 VDD sg13_lv_pmos w={CP_P_W} l={CP_P_L} ng=1 m={CP_P_M}
XM10 net4 UP VDD VDD sg13_lv_pmos w={CP_P_W} l={CP_P_L} ng=1 m={CP_P_M}
XC1 net5 GND cparasitic C='C_CP'
XR1 Ibias Vbp sub! rsil w=0.5e-6 l=0.5e-6 m=1 b=0
XM11 VDD net5 CTRL GND sg13_lv_nmos w=100u l=0.5u ng=20 m=1
XR2 GND CTRL sub! rsil w=0.5e-6 l=0.5e-4 m=1 b=0
XR3 net6 net5 sub! rsil w=0.5e-6 l=1e-5 m=1 b=0
.ends


* expanding   symbol:  /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/phase-freq-detector/PFD_std.sym # of
*+ pins=6
** sym_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/phase-freq-detector/PFD_std.sym
** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/phase-freq-detector/PFD_std.sch
.subckt PFD_std VDD UP F_REF F_VCO DN GND
*.opin UP
*.ipin F_REF
*.ipin VDD
*.ipin GND
*.opin DN
*.ipin F_VCO
x1 net1 net2 F_REF VDD RST_N VDD GND sg13g2_dfrbp_2
x2 DN net3 F_VCO VDD RST_N VDD GND sg13g2_dfrbp_2
x3 RST_N net1 DN VDD GND sg13g2_nand2_2
x4 UP net1 VDD GND sg13g2_inv_2
.ends


* expanding   symbol:  /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/top-pll/FD/Freq_Div_std.sym # of
*+ pins=2
** sym_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/top-pll/FD/Freq_Div_std.sym
** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/top-pll/FD/Freq_Div_std.sch
.subckt Freq_Div_std F_IN F_OUT
*.opin F_OUT
*.ipin F_IN
x6 net3 net1 F_IN net1 VDD VDD GND sg13g2_dfrbp_1
x5 net4 net2 net3 net2 VDD VDD GND sg13g2_dfrbp_2
x7 net6 net5 net4 net5 VDD VDD GND sg13g2_dfrbp_2
x8 F_OUT net7 net6 net7 VDD VDD GND sg13g2_dfrbp_2
.ends

.GLOBAL GND
.GLOBAL VDD
.end
