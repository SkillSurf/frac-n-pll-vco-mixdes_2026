* Extracted by KLayout with SG13G2 LVS runset on : 13/07/2025 18:41

.SUBCKT TOP
X$1 13 12 9 1 12 pmos$1
X$2 13 8 9 1 8 pmos$2
X$3 6 11 6 9 1 8 8 pmos
X$4 8 7 1 10 nmos$1
X$5 10 2 1 6 nmos$2
X$6 13 11 1 rppd$1
X$7 2 3 1 rppd$1
X$8 8 3 1 6 nmos$2
X$9 6 2 1 6 nmos$2
X$10 6 2 1 4 nmos$1
X$11 7 2 1 5 nmos$1
X$12 13 8 9 1 5 pmos$1
X$13 12 10 9 1 10 pmos$1
X$14 13 10 9 1 5 pmos$1
.ENDS TOP

.SUBCKT rppd$1 1 2 3
R$1 1 2 rppd w=1u l=12u ps=0 b=0 m=1
.ENDS rppd$1

.SUBCKT nmos$2 1 2 3 4
M$1 1 4 2 3 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
.ENDS nmos$2

.SUBCKT nmos$1 1 2 3 4
M$1 1 4 2 3 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
.ENDS nmos$1

.SUBCKT pmos 1 2 3 4 5 6 7
M$1 1 6 2 4 sg13_lv_pmos L=1u W=2u AS=0.68p AD=0.38p PS=4.68u PD=2.38u
M$2 2 7 3 4 sg13_lv_pmos L=1u W=2u AS=0.38p AD=0.68p PS=2.38u PD=4.68u
.ENDS pmos

.SUBCKT pmos$2 1 2 3 4 5
M$1 1 5 2 3 sg13_lv_pmos L=1u W=2u AS=0.68p AD=0.68p PS=4.68u PD=4.68u
.ENDS pmos$2

.SUBCKT pmos$1 1 2 3 4 5
M$1 1 5 2 3 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
.ENDS pmos$1
