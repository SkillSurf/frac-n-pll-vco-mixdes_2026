** sch_path: /home/mmhnbm/frac-n-pll-vco-smacd_2026/schematic/blocks/dsm/xschem/dsm_with_mdiv_tb.sch
**.subckt dsm_with_mdiv_tb
V1 freq_in GND PULSE(0 1.8 0 10ns 10ns 50ns 100ns)
A2 [ en ] [ net2 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=1.2
A3 [ sdata ] [ net3 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=1.2
A4 [ sclk ] [ net4 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=1.2
A5 [ rst ] [ net5 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=1.2
A6 [ freq_in ] [ net6 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=1.2
* noconn rst
* noconn sclk
* noconn sdata
* noconn en
A10 [ net1 ] [ freq_out ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
adut [ net6 net5 net4 net3 net2 ] [ net1 ] null dut
.model dut d_cosim simulation=./../dsm_and_freq_divider.so
**** begin user architecture code



* ngspice commands
.save v(dout) v(sdata) v(sclk) v(en) v(rst) v(dsm_clk) v(freq_in) v(freq_out)
.control
  tran 0.5n 1m
  remzerovec
  write test.raw
.endc

* to generate following file copy stimuli.test
* to the simulation directory and run simulation -> Utile Stimuli Editor (GUI),
* and press 'Translate'
.include stimuli_test.cir


**** end user architecture code
**.ends
.GLOBAL GND
.end
