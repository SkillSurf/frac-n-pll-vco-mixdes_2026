.subckt IHP_4nH_Inductor 1 2
Vam1 1 n2 dc 0
Rport1 n2 0 50
Vam2 2 n4 dc 0
Rport2 n4 0 50

Fi1 0 ni1 Vam1 50
Gi1 0 ni1 1 0 1
Rt1 ni1 0 1
Fi2 0 ni2 Vam2 50
Gi2 0 ni2 2 0 1
Rt2 ni2 0 1

Ca1 ns1 0 1e-012
Ra1 ns1 0 131834.068078
Ca2 ns2 0 1e-012
Ra2 ns2 0 735.819681122
Ca3 ns3 0 1e-012
Ca4 ns4 0 1e-012
Ra3 ns3 0 186.359484923
Ra4 ns4 0 186.359484923
Ga3 ns3 0 ns4 0 -0.00231880636624
Ga4 ns4 0 ns3 0 0.00231880636624
Ca5 ns5 0 1e-012
Ra5 ns5 0 141.613068254
Ca6 ns6 0 1e-012
Ra6 ns6 0 29.4273648628
Ca7 ns7 0 1e-012
Ca8 ns8 0 1e-012
Ra7 ns7 0 8.35389829092
Ra8 ns8 0 8.35389829092
Ga7 ns7 0 ns8 0 -0.17749287689
Ga8 ns8 0 ns7 0 0.17749287689
Ca9 ns9 0 1e-012
Ra9 ns9 0 3.07433189927
Ca10 ns10 0 1e-012
Ra10 ns10 0 131834.068078
Ca11 ns11 0 1e-012
Ra11 ns11 0 735.819681122
Ca12 ns12 0 1e-012
Ca13 ns13 0 1e-012
Ra12 ns12 0 186.359484923
Ra13 ns13 0 186.359484923
Ga12 ns12 0 ns13 0 -0.00231880636624
Ga13 ns13 0 ns12 0 0.00231880636624
Ca14 ns14 0 1e-012
Ra14 ns14 0 141.613068254
Ca15 ns15 0 1e-012
Ra15 ns15 0 29.4273648628
Ca16 ns16 0 1e-012
Ca17 ns17 0 1e-012
Ra16 ns16 0 8.35389829092
Ra17 ns17 0 8.35389829092
Ga16 ns16 0 ns17 0 -0.17749287689
Ga17 ns17 0 ns16 0 0.17749287689
Ca18 ns18 0 1e-012
Ra18 ns18 0 3.07433189927

Gb1_1 ns1 0 ni1 0 7.58529274395e-006
Gb2_1 ns2 0 ni1 0 0.00135902861211
Gb3_1 ns3 0 ni1 0 0.00636800260357
Gb5_1 ns5 0 ni1 0 0.00706149518775
Gb6_1 ns6 0 ni1 0 0.0339819757788
Gb7_1 ns7 0 ni1 0 0.25822394612
Gb9_1 ns9 0 ni1 0 0.32527392382
Gb10_2 ns10 0 ni2 0 7.58529274395e-006
Gb11_2 ns11 0 ni2 0 0.00135902861211
Gb12_2 ns12 0 ni2 0 0.00636800260357
Gb14_2 ns14 0 ni2 0 0.00706149518775
Gb15_2 ns15 0 ni2 0 0.0339819757788
Gb16_2 ns16 0 ni2 0 0.25822394612
Gb18_2 ns18 0 ni2 0 0.32527392382

Gc1_1 0 n2 ns1 0 2.84507160964e-005
Gc1_2 0 n2 ns2 0 -0.000166153915314
Gc1_3 0 n2 ns3 0 -0.000263626276308
Gc1_4 0 n2 ns4 0 -1.97468499264e-005
Gc1_5 0 n2 ns5 0 0.000589105007869
Gc1_6 0 n2 ns6 0 0.0316346578419
Gc1_7 0 n2 ns7 0 0.0365168086279
Gc1_8 0 n2 ns8 0 -0.00235594459174
Gc1_9 0 n2 ns9 0 -0.0695812178423
Gc1_10 0 n2 ns10 0 -2.8091743964e-005
Gc1_11 0 n2 ns11 0 -0.000235604054074
Gc1_12 0 n2 ns12 0 0.000403582669599
Gc1_13 0 n2 ns13 0 9.09461127e-005
Gc1_14 0 n2 ns14 0 -0.000951296496322
Gc1_15 0 n2 ns15 0 -0.0316664072649
Gc1_16 0 n2 ns16 0 -0.03768425623
Gc1_17 0 n2 ns17 0 0.00504639696586
Gc1_18 0 n2 ns18 0 0.0451786493797
Gd1_1 0 n2 ni1 0 -0.0105028683359
Gd1_2 0 n2 ni2 0 0.00193597863844
Gc2_1 0 n4 ns1 0 -2.80917439638e-005
Gc2_2 0 n4 ns2 0 -0.000235604054075
Gc2_3 0 n4 ns3 0 0.000403582669594
Gc2_4 0 n4 ns4 0 9.09461126972e-005
Gc2_5 0 n4 ns5 0 -0.000951296496319
Gc2_6 0 n4 ns6 0 -0.0316664072649
Gc2_7 0 n4 ns7 0 -0.03768425623
Gc2_8 0 n4 ns8 0 0.00504639696583
Gc2_9 0 n4 ns9 0 0.0451786493796
Gc2_10 0 n4 ns10 0 2.85337921315e-005
Gc2_11 0 n4 ns11 0 -0.000168536641816
Gc2_12 0 n4 ns12 0 -0.000272282905638
Gc2_13 0 n4 ns13 0 -2.42792134581e-005
Gc2_14 0 n4 ns14 0 0.000591575130422
Gc2_15 0 n4 ns15 0 0.0316267338258
Gc2_16 0 n4 ns16 0 0.0354660552526
Gc2_17 0 n4 ns17 0 -0.00282616402358
Gc2_18 0 n4 ns18 0 -0.0703910464608
Gd2_1 0 n4 ni1 0 0.00193597863841
Gd2_2 0 n4 ni2 0 -0.0115657051542
.ends
