** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/top-pll/Frequency_Divider_tb.sch
**.subckt Frequency_Divider_tb
V1 VDD GND 1.2
Vfref F_REF GND 0 pulse(0 1.2 0p 100p 100p 200p 400p)
x1 F_REF F_OUT Freq_Div_std
**** begin user architecture code



.model freq_div freq_div
*.include tb_CP.save
.param RAW_TEMP = agauss(40, 30, 1)
.param TEMPGAUSS = max(20, min(RAW_TEMP, 80))
.option temp = 'TEMPGAUSS'
.param VDDGAUSS = agauss(1.2, 0.05, 1)

.param VDD = 'VDDGAUSS'
* analysis

.control
pre_osdi /foss/designs/PLL_IHP_PDK/src/freq_div.osdi
save all
write Frequency_divider_tb.raw
set appendwrite
let i = 0
dowhile i < 1


  tran 10p 200n uic
  write tb_Frequency_Divisder.raw
  linearize
  fft v(F_REF) v(F_OUT)
  write tb_Frequency_Divisder.raw
  let i = i + 1
end
*quit 0
.endc





.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ_stat
.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice
.global VDD GND


**** end user architecture code
**.ends

* expanding   symbol:  Freq_Div_std.sym # of pins=2
** sym_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/top-pll/Freq_Div_std.sym
** sch_path: /foss/designs/iic_osic_tools/frac-n-pll-vco-unic_cass/schematic/blocks/top-pll/Freq_Div_std.sch
.subckt Freq_Div_std F_IN F_OUT
*.opin F_OUT
*.ipin F_IN
x6 net3 net1 F_IN net1 VDD VDD GND sg13g2_dfrbp_1
x5 net4 net2 net3 net2 VDD VDD GND sg13g2_dfrbp_2
x7 net6 net5 net4 net5 VDD VDD GND sg13g2_dfrbp_2
x8 F_OUT net7 net6 net7 VDD VDD GND sg13g2_dfrbp_2
.ends

.GLOBAL GND
.GLOBAL VDD
.end
